module game_logic_top();

// 

endmodule