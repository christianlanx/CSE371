module fifo_buffer() 